module top_module( input in, output out );

    // veriog has bit-wise NOT (~) and logical NOT (!)
    assign out = ~in;
    
endmodule
